-- Garfield_system.vhd

-- Generated using ACDS version 16.0 222

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Garfield_system is
	port (
		clk_clk                                          : in    std_logic                     := '0';             --                                       clk.clk
		clk_1_fpga_clock_clk                             : in    std_logic                     := '0';             --                          clk_1_fpga_clock.clk
		clk_1_fpga_reset_reset_n                         : in    std_logic                     := '0';             --                          clk_1_fpga_reset.reset_n
		garfield_general_io_external_connection_export   : out   std_logic_vector(7 downto 0);                     --   garfield_general_io_external_connection.export
		garfield_lighting_led_external_connection_export : out   std_logic_vector(3 downto 0);                     -- garfield_lighting_led_external_connection.export
		hps_0_f2h_cold_reset_req_reset_n                 : in    std_logic                     := '0';             --                  hps_0_f2h_cold_reset_req.reset_n
		hps_0_f2h_debug_reset_req_reset_n                : in    std_logic                     := '0';             --                 hps_0_f2h_debug_reset_req.reset_n
		hps_0_f2h_stm_hw_events_stm_hwevents             : in    std_logic_vector(27 downto 0) := (others => '0'); --                   hps_0_f2h_stm_hw_events.stm_hwevents
		hps_0_f2h_warm_reset_req_reset_n                 : in    std_logic                     := '0';             --                  hps_0_f2h_warm_reset_req.reset_n
		hps_0_h2f_reset_reset_n                          : out   std_logic;                                        --                           hps_0_h2f_reset.reset_n
		hps_0_hps_io_hps_io_emac1_inst_TX_CLK            : out   std_logic;                                        --                              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		hps_0_hps_io_hps_io_emac1_inst_TXD0              : out   std_logic;                                        --                                          .hps_io_emac1_inst_TXD0
		hps_0_hps_io_hps_io_emac1_inst_TXD1              : out   std_logic;                                        --                                          .hps_io_emac1_inst_TXD1
		hps_0_hps_io_hps_io_emac1_inst_TXD2              : out   std_logic;                                        --                                          .hps_io_emac1_inst_TXD2
		hps_0_hps_io_hps_io_emac1_inst_TXD3              : out   std_logic;                                        --                                          .hps_io_emac1_inst_TXD3
		hps_0_hps_io_hps_io_emac1_inst_RXD0              : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RXD0
		hps_0_hps_io_hps_io_emac1_inst_MDIO              : inout std_logic                     := '0';             --                                          .hps_io_emac1_inst_MDIO
		hps_0_hps_io_hps_io_emac1_inst_MDC               : out   std_logic;                                        --                                          .hps_io_emac1_inst_MDC
		hps_0_hps_io_hps_io_emac1_inst_RX_CTL            : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RX_CTL
		hps_0_hps_io_hps_io_emac1_inst_TX_CTL            : out   std_logic;                                        --                                          .hps_io_emac1_inst_TX_CTL
		hps_0_hps_io_hps_io_emac1_inst_RX_CLK            : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RX_CLK
		hps_0_hps_io_hps_io_emac1_inst_RXD1              : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RXD1
		hps_0_hps_io_hps_io_emac1_inst_RXD2              : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RXD2
		hps_0_hps_io_hps_io_emac1_inst_RXD3              : in    std_logic                     := '0';             --                                          .hps_io_emac1_inst_RXD3
		hps_0_hps_io_hps_io_sdio_inst_CMD                : inout std_logic                     := '0';             --                                          .hps_io_sdio_inst_CMD
		hps_0_hps_io_hps_io_sdio_inst_D0                 : inout std_logic                     := '0';             --                                          .hps_io_sdio_inst_D0
		hps_0_hps_io_hps_io_sdio_inst_D1                 : inout std_logic                     := '0';             --                                          .hps_io_sdio_inst_D1
		hps_0_hps_io_hps_io_sdio_inst_CLK                : out   std_logic;                                        --                                          .hps_io_sdio_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_D2                 : inout std_logic                     := '0';             --                                          .hps_io_sdio_inst_D2
		hps_0_hps_io_hps_io_sdio_inst_D3                 : inout std_logic                     := '0';             --                                          .hps_io_sdio_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D0                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D0
		hps_0_hps_io_hps_io_usb1_inst_D1                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D1
		hps_0_hps_io_hps_io_usb1_inst_D2                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D2
		hps_0_hps_io_hps_io_usb1_inst_D3                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D4                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D4
		hps_0_hps_io_hps_io_usb1_inst_D5                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D5
		hps_0_hps_io_hps_io_usb1_inst_D6                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D6
		hps_0_hps_io_hps_io_usb1_inst_D7                 : inout std_logic                     := '0';             --                                          .hps_io_usb1_inst_D7
		hps_0_hps_io_hps_io_usb1_inst_CLK                : in    std_logic                     := '0';             --                                          .hps_io_usb1_inst_CLK
		hps_0_hps_io_hps_io_usb1_inst_STP                : out   std_logic;                                        --                                          .hps_io_usb1_inst_STP
		hps_0_hps_io_hps_io_usb1_inst_DIR                : in    std_logic                     := '0';             --                                          .hps_io_usb1_inst_DIR
		hps_0_hps_io_hps_io_usb1_inst_NXT                : in    std_logic                     := '0';             --                                          .hps_io_usb1_inst_NXT
		hps_0_hps_io_hps_io_spim1_inst_CLK               : out   std_logic;                                        --                                          .hps_io_spim1_inst_CLK
		hps_0_hps_io_hps_io_spim1_inst_MOSI              : out   std_logic;                                        --                                          .hps_io_spim1_inst_MOSI
		hps_0_hps_io_hps_io_spim1_inst_MISO              : in    std_logic                     := '0';             --                                          .hps_io_spim1_inst_MISO
		hps_0_hps_io_hps_io_spim1_inst_SS0               : out   std_logic;                                        --                                          .hps_io_spim1_inst_SS0
		hps_0_hps_io_hps_io_uart0_inst_RX                : in    std_logic                     := '0';             --                                          .hps_io_uart0_inst_RX
		hps_0_hps_io_hps_io_uart0_inst_TX                : out   std_logic;                                        --                                          .hps_io_uart0_inst_TX
		hps_0_hps_io_hps_io_i2c0_inst_SDA                : inout std_logic                     := '0';             --                                          .hps_io_i2c0_inst_SDA
		hps_0_hps_io_hps_io_i2c0_inst_SCL                : inout std_logic                     := '0';             --                                          .hps_io_i2c0_inst_SCL
		hps_0_hps_io_hps_io_i2c1_inst_SDA                : inout std_logic                     := '0';             --                                          .hps_io_i2c1_inst_SDA
		hps_0_hps_io_hps_io_i2c1_inst_SCL                : inout std_logic                     := '0';             --                                          .hps_io_i2c1_inst_SCL
		hps_0_hps_io_hps_io_gpio_inst_GPIO09             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO09
		hps_0_hps_io_hps_io_gpio_inst_GPIO35             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO35
		hps_0_hps_io_hps_io_gpio_inst_GPIO40             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO40
		hps_0_hps_io_hps_io_gpio_inst_GPIO53             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO53
		hps_0_hps_io_hps_io_gpio_inst_GPIO54             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO54
		hps_0_hps_io_hps_io_gpio_inst_GPIO61             : inout std_logic                     := '0';             --                                          .hps_io_gpio_inst_GPIO61
		i2c_0_external_connection_scl_pad_io             : inout std_logic                     := '0';             --                 i2c_0_external_connection.scl_pad_io
		i2c_0_external_connection_sda_pad_io             : inout std_logic                     := '0';             --                                          .sda_pad_io
		memory_mem_a                                     : out   std_logic_vector(14 downto 0);                    --                                    memory.mem_a
		memory_mem_ba                                    : out   std_logic_vector(2 downto 0);                     --                                          .mem_ba
		memory_mem_ck                                    : out   std_logic;                                        --                                          .mem_ck
		memory_mem_ck_n                                  : out   std_logic;                                        --                                          .mem_ck_n
		memory_mem_cke                                   : out   std_logic;                                        --                                          .mem_cke
		memory_mem_cs_n                                  : out   std_logic;                                        --                                          .mem_cs_n
		memory_mem_ras_n                                 : out   std_logic;                                        --                                          .mem_ras_n
		memory_mem_cas_n                                 : out   std_logic;                                        --                                          .mem_cas_n
		memory_mem_we_n                                  : out   std_logic;                                        --                                          .mem_we_n
		memory_mem_reset_n                               : out   std_logic;                                        --                                          .mem_reset_n
		memory_mem_dq                                    : inout std_logic_vector(31 downto 0) := (others => '0'); --                                          .mem_dq
		memory_mem_dqs                                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                          .mem_dqs
		memory_mem_dqs_n                                 : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                          .mem_dqs_n
		memory_mem_odt                                   : out   std_logic;                                        --                                          .mem_odt
		memory_mem_dm                                    : out   std_logic_vector(3 downto 0);                     --                                          .mem_dm
		memory_oct_rzqin                                 : in    std_logic                     := '0';             --                                          .oct_rzqin
		onboard_button_external_connection_export        : in    std_logic_vector(1 downto 0)  := (others => '0'); --        onboard_button_external_connection.export
		onboard_dipsw_external_connection_export         : in    std_logic_vector(3 downto 0)  := (others => '0'); --         onboard_dipsw_external_connection.export
		onboard_led_external_connection_export           : out   std_logic_vector(7 downto 0);                     --           onboard_led_external_connection.export
		reset_reset_n                                    : in    std_logic                     := '0';             --                                     reset.reset_n
		spi_0_external_connection_MISO                   : in    std_logic                     := '0';             --                 spi_0_external_connection.MISO
		spi_0_external_connection_MOSI                   : out   std_logic;                                        --                                          .MOSI
		spi_0_external_connection_SCLK                   : out   std_logic;                                        --                                          .SCLK
		spi_0_external_connection_SS_n                   : out   std_logic_vector(2 downto 0)                      --                                          .SS_n
	);
end entity Garfield_system;

architecture rtl of Garfield_system is
	component Garfield_system_Garfield_GPIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Garfield_system_Garfield_GPIO;

	component Garfield_system_Garfield_lighting is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component Garfield_system_Garfield_lighting;

	component Garfield_system_Onboard_Button is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component Garfield_system_Onboard_Button;

	component Garfield_system_Onboard_DipSW is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component Garfield_system_Onboard_DipSW;

	component Garfield_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_cold_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			f2h_dbg_rst_req_n        : in    std_logic                      := 'X';             -- reset_n
			f2h_warm_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0)  := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component Garfield_system_hps_0;

	component i2c_opencores is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component Garfield_system_jtag_uart_nios2 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Garfield_system_jtag_uart_nios2;

	component Garfield_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(22 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Garfield_system_nios2_gen2_0;

	component Garfield_system_onchip_memory2_nios2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component Garfield_system_onchip_memory2_nios2;

	component Garfield_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Garfield_system_pll_0;

	component Garfield_system_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(2 downto 0)                      -- export
		);
	end component Garfield_system_spi_0;

	component Garfield_system_sysid_fpga is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Garfield_system_sysid_fpga;

	component Garfield_system_timer_0_nios2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Garfield_system_timer_0_nios2;

	component Garfield_system_mm_interconnect_0 is
		port (
			pll_0_outclk0_clk                              : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			Garfield_GPIO_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			Garfield_GPIO_s1_write                         : out std_logic;                                        -- write
			Garfield_GPIO_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Garfield_GPIO_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			Garfield_GPIO_s1_chipselect                    : out std_logic;                                        -- chipselect
			Garfield_lighting_s1_address                   : out std_logic_vector(1 downto 0);                     -- address
			Garfield_lighting_s1_write                     : out std_logic;                                        -- write
			Garfield_lighting_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Garfield_lighting_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			Garfield_lighting_s1_chipselect                : out std_logic;                                        -- chipselect
			i2c_opencores_0_avalon_slave_0_address         : out std_logic_vector(2 downto 0);                     -- address
			i2c_opencores_0_avalon_slave_0_write           : out std_logic;                                        -- write
			i2c_opencores_0_avalon_slave_0_readdata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_opencores_0_avalon_slave_0_writedata       : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_opencores_0_avalon_slave_0_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect      : out std_logic;                                        -- chipselect
			jtag_uart_nios2_avalon_jtag_slave_address      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_nios2_avalon_jtag_slave_write        : out std_logic;                                        -- write
			jtag_uart_nios2_avalon_jtag_slave_read         : out std_logic;                                        -- read
			jtag_uart_nios2_avalon_jtag_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_nios2_avalon_jtag_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_nios2_avalon_jtag_slave_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_nios2_avalon_jtag_slave_chipselect   : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			Onboard_Button_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			Onboard_Button_s1_write                        : out std_logic;                                        -- write
			Onboard_Button_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onboard_Button_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			Onboard_Button_s1_chipselect                   : out std_logic;                                        -- chipselect
			Onboard_DipSW_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			Onboard_DipSW_s1_write                         : out std_logic;                                        -- write
			Onboard_DipSW_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onboard_DipSW_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			Onboard_DipSW_s1_chipselect                    : out std_logic;                                        -- chipselect
			Onboard_LED_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			Onboard_LED_s1_write                           : out std_logic;                                        -- write
			Onboard_LED_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onboard_LED_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Onboard_LED_s1_chipselect                      : out std_logic;                                        -- chipselect
			onchip_memory2_nios2_s1_address                : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_nios2_s1_write                  : out std_logic;                                        -- write
			onchip_memory2_nios2_s1_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_nios2_s1_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_nios2_s1_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_nios2_s1_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory2_nios2_s1_clken                  : out std_logic;                                        -- clken
			spi_0_spi_control_port_address                 : out std_logic_vector(2 downto 0);                     -- address
			spi_0_spi_control_port_write                   : out std_logic;                                        -- write
			spi_0_spi_control_port_read                    : out std_logic;                                        -- read
			spi_0_spi_control_port_readdata                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_0_spi_control_port_writedata               : out std_logic_vector(15 downto 0);                    -- writedata
			spi_0_spi_control_port_chipselect              : out std_logic;                                        -- chipselect
			sysid_fpga_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_fpga_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_nios2_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			timer_0_nios2_s1_write                         : out std_logic;                                        -- write
			timer_0_nios2_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_nios2_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_nios2_s1_chipselect                    : out std_logic                                         -- chipselect
		);
	end component Garfield_system_mm_interconnect_0;

	component Garfield_system_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Garfield_system_irq_mapper;

	component Garfield_system_irq_mapper_002 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Garfield_system_irq_mapper_002;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal pll_0_outclk0_clk                                                   : std_logic;                     -- pll_0:outclk_0 -> [Garfield_GPIO:clk, Garfield_lighting:clk, Onboard_Button:clk, Onboard_DipSW:clk, Onboard_LED:clk, i2c_opencores_0:wb_clk_i, irq_mapper_002:clk, jtag_uart_nios2:clk, mm_interconnect_0:pll_0_outclk0_clk, nios2_gen2_0:clk, onchip_memory2_nios2:clk, rst_controller:clk, spi_0:clk, sysid_fpga:clock, timer_0_nios2:clk]
	signal nios2_gen2_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                    : std_logic_vector(22 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                       : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                      : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                             : std_logic_vector(18 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_chipselect -> jtag_uart_nios2:av_chipselect
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_nios2:av_readdata -> mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_nios2:av_waitrequest -> mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_address -> jtag_uart_nios2:av_address
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_nios2_avalon_jtag_slave_writedata -> jtag_uart_nios2:av_writedata
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect         : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata           : std_logic_vector(7 downto 0);  -- i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	signal i2c_opencores_0_avalon_slave_0_waitrequest                          : std_logic;                     -- i2c_opencores_0:wb_ack_o -> i2c_opencores_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write              : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	signal mm_interconnect_0_sysid_fpga_control_slave_readdata                 : std_logic_vector(31 downto 0); -- sysid_fpga:readdata -> mm_interconnect_0:sysid_fpga_control_slave_readdata
	signal mm_interconnect_0_sysid_fpga_control_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_fpga_control_slave_address -> sysid_fpga:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest          : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_nios2_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_nios2_s1_chipselect -> onchip_memory2_nios2:chipselect
	signal mm_interconnect_0_onchip_memory2_nios2_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_nios2:readdata -> mm_interconnect_0:onchip_memory2_nios2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_nios2_s1_address                   : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_nios2_s1_address -> onchip_memory2_nios2:address
	signal mm_interconnect_0_onchip_memory2_nios2_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_nios2_s1_byteenable -> onchip_memory2_nios2:byteenable
	signal mm_interconnect_0_onchip_memory2_nios2_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_nios2_s1_write -> onchip_memory2_nios2:write
	signal mm_interconnect_0_onchip_memory2_nios2_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_nios2_s1_writedata -> onchip_memory2_nios2:writedata
	signal mm_interconnect_0_onchip_memory2_nios2_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_nios2_s1_clken -> onchip_memory2_nios2:clken
	signal mm_interconnect_0_onboard_led_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:Onboard_LED_s1_chipselect -> Onboard_LED:chipselect
	signal mm_interconnect_0_onboard_led_s1_readdata                           : std_logic_vector(31 downto 0); -- Onboard_LED:readdata -> mm_interconnect_0:Onboard_LED_s1_readdata
	signal mm_interconnect_0_onboard_led_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Onboard_LED_s1_address -> Onboard_LED:address
	signal mm_interconnect_0_onboard_led_s1_write                              : std_logic;                     -- mm_interconnect_0:Onboard_LED_s1_write -> mm_interconnect_0_onboard_led_s1_write:in
	signal mm_interconnect_0_onboard_led_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onboard_LED_s1_writedata -> Onboard_LED:writedata
	signal mm_interconnect_0_onboard_button_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:Onboard_Button_s1_chipselect -> Onboard_Button:chipselect
	signal mm_interconnect_0_onboard_button_s1_readdata                        : std_logic_vector(31 downto 0); -- Onboard_Button:readdata -> mm_interconnect_0:Onboard_Button_s1_readdata
	signal mm_interconnect_0_onboard_button_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Onboard_Button_s1_address -> Onboard_Button:address
	signal mm_interconnect_0_onboard_button_s1_write                           : std_logic;                     -- mm_interconnect_0:Onboard_Button_s1_write -> mm_interconnect_0_onboard_button_s1_write:in
	signal mm_interconnect_0_onboard_button_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onboard_Button_s1_writedata -> Onboard_Button:writedata
	signal mm_interconnect_0_onboard_dipsw_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Onboard_DipSW_s1_chipselect -> Onboard_DipSW:chipselect
	signal mm_interconnect_0_onboard_dipsw_s1_readdata                         : std_logic_vector(31 downto 0); -- Onboard_DipSW:readdata -> mm_interconnect_0:Onboard_DipSW_s1_readdata
	signal mm_interconnect_0_onboard_dipsw_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Onboard_DipSW_s1_address -> Onboard_DipSW:address
	signal mm_interconnect_0_onboard_dipsw_s1_write                            : std_logic;                     -- mm_interconnect_0:Onboard_DipSW_s1_write -> mm_interconnect_0_onboard_dipsw_s1_write:in
	signal mm_interconnect_0_onboard_dipsw_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onboard_DipSW_s1_writedata -> Onboard_DipSW:writedata
	signal mm_interconnect_0_timer_0_nios2_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:timer_0_nios2_s1_chipselect -> timer_0_nios2:chipselect
	signal mm_interconnect_0_timer_0_nios2_s1_readdata                         : std_logic_vector(15 downto 0); -- timer_0_nios2:readdata -> mm_interconnect_0:timer_0_nios2_s1_readdata
	signal mm_interconnect_0_timer_0_nios2_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_nios2_s1_address -> timer_0_nios2:address
	signal mm_interconnect_0_timer_0_nios2_s1_write                            : std_logic;                     -- mm_interconnect_0:timer_0_nios2_s1_write -> mm_interconnect_0_timer_0_nios2_s1_write:in
	signal mm_interconnect_0_timer_0_nios2_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_nios2_s1_writedata -> timer_0_nios2:writedata
	signal mm_interconnect_0_garfield_lighting_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:Garfield_lighting_s1_chipselect -> Garfield_lighting:chipselect
	signal mm_interconnect_0_garfield_lighting_s1_readdata                     : std_logic_vector(31 downto 0); -- Garfield_lighting:readdata -> mm_interconnect_0:Garfield_lighting_s1_readdata
	signal mm_interconnect_0_garfield_lighting_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Garfield_lighting_s1_address -> Garfield_lighting:address
	signal mm_interconnect_0_garfield_lighting_s1_write                        : std_logic;                     -- mm_interconnect_0:Garfield_lighting_s1_write -> mm_interconnect_0_garfield_lighting_s1_write:in
	signal mm_interconnect_0_garfield_lighting_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:Garfield_lighting_s1_writedata -> Garfield_lighting:writedata
	signal mm_interconnect_0_garfield_gpio_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:Garfield_GPIO_s1_chipselect -> Garfield_GPIO:chipselect
	signal mm_interconnect_0_garfield_gpio_s1_readdata                         : std_logic_vector(31 downto 0); -- Garfield_GPIO:readdata -> mm_interconnect_0:Garfield_GPIO_s1_readdata
	signal mm_interconnect_0_garfield_gpio_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Garfield_GPIO_s1_address -> Garfield_GPIO:address
	signal mm_interconnect_0_garfield_gpio_s1_write                            : std_logic;                     -- mm_interconnect_0:Garfield_GPIO_s1_write -> mm_interconnect_0_garfield_gpio_s1_write:in
	signal mm_interconnect_0_garfield_gpio_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:Garfield_GPIO_s1_writedata -> Garfield_GPIO:writedata
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect                 : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata                   : std_logic_vector(15 downto 0); -- spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                       : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write                      : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	signal hps_0_f2h_irq0_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal irq_mapper_002_receiver0_irq                                        : std_logic;                     -- i2c_opencores_0:wb_inta_o -> irq_mapper_002:receiver0_irq
	signal irq_mapper_002_receiver1_irq                                        : std_logic;                     -- jtag_uart_nios2:av_irq -> irq_mapper_002:receiver1_irq
	signal irq_mapper_002_receiver2_irq                                        : std_logic;                     -- timer_0_nios2:irq -> irq_mapper_002:receiver2_irq
	signal irq_mapper_002_receiver3_irq                                        : std_logic;                     -- spi_0:irq -> irq_mapper_002:receiver3_irq
	signal nios2_gen2_0_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [i2c_opencores_0:wb_rst_i, irq_mapper_002:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_nios2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_nios2:reset_req, rst_translator:reset_req_in]
	signal clk_1_fpga_reset_reset_n_ports_inv                                  : std_logic;                     -- clk_1_fpga_reset_reset_n:inv -> [pll_0:rst, rst_controller:reset_in0]
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read:inv -> jtag_uart_nios2:av_read_n
	signal mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write:inv -> jtag_uart_nios2:av_write_n
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv                : std_logic;                     -- i2c_opencores_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_onboard_led_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_onboard_led_s1_write:inv -> Onboard_LED:write_n
	signal mm_interconnect_0_onboard_button_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_onboard_button_s1_write:inv -> Onboard_Button:write_n
	signal mm_interconnect_0_onboard_dipsw_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_onboard_dipsw_s1_write:inv -> Onboard_DipSW:write_n
	signal mm_interconnect_0_timer_0_nios2_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_timer_0_nios2_s1_write:inv -> timer_0_nios2:write_n
	signal mm_interconnect_0_garfield_lighting_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_garfield_lighting_s1_write:inv -> Garfield_lighting:write_n
	signal mm_interconnect_0_garfield_gpio_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_garfield_gpio_s1_write:inv -> Garfield_GPIO:write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv             : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> spi_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv            : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> spi_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Garfield_GPIO:reset_n, Garfield_lighting:reset_n, Onboard_Button:reset_n, Onboard_DipSW:reset_n, Onboard_LED:reset_n, jtag_uart_nios2:rst_n, nios2_gen2_0:reset_n, spi_0:reset_n, sysid_fpga:reset_n, timer_0_nios2:reset_n]

begin

	garfield_gpio : component Garfield_system_Garfield_GPIO
		port map (
			clk        => pll_0_outclk0_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_garfield_gpio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_garfield_gpio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_garfield_gpio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_garfield_gpio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_garfield_gpio_s1_readdata,        --                    .readdata
			out_port   => garfield_general_io_external_connection_export      -- external_connection.export
		);

	garfield_lighting : component Garfield_system_Garfield_lighting
		port map (
			clk        => pll_0_outclk0_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => mm_interconnect_0_garfield_lighting_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_garfield_lighting_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_garfield_lighting_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_garfield_lighting_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_garfield_lighting_s1_readdata,        --                    .readdata
			out_port   => garfield_lighting_led_external_connection_export        -- external_connection.export
		);

	onboard_button : component Garfield_system_Onboard_Button
		port map (
			clk        => pll_0_outclk0_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_onboard_button_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_onboard_button_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_onboard_button_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_onboard_button_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_onboard_button_s1_readdata,        --                    .readdata
			in_port    => onboard_button_external_connection_export            -- external_connection.export
		);

	onboard_dipsw : component Garfield_system_Onboard_DipSW
		port map (
			clk        => pll_0_outclk0_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_onboard_dipsw_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_onboard_dipsw_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_onboard_dipsw_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_onboard_dipsw_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_onboard_dipsw_s1_readdata,        --                    .readdata
			in_port    => onboard_dipsw_external_connection_export            -- external_connection.export
		);

	onboard_led : component Garfield_system_Garfield_GPIO
		port map (
			clk        => pll_0_outclk0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_onboard_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_onboard_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_onboard_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_onboard_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_onboard_led_s1_readdata,        --                    .readdata
			out_port   => onboard_led_external_connection_export            -- external_connection.export
		);

	hps_0 : component Garfield_system_hps_0
		generic map (
			F2S_Width => 3,
			S2F_Width => 2
		)
		port map (
			f2h_cold_rst_req_n       => hps_0_f2h_cold_reset_req_reset_n,      --  f2h_cold_reset_req.reset_n
			f2h_dbg_rst_req_n        => hps_0_f2h_debug_reset_req_reset_n,     -- f2h_debug_reset_req.reset_n
			f2h_warm_rst_req_n       => hps_0_f2h_warm_reset_req_reset_n,      --  f2h_warm_reset_req.reset_n
			f2h_stm_hwevents         => hps_0_f2h_stm_hw_events_stm_hwevents,  --   f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                          --              memory.mem_a
			mem_ba                   => memory_mem_ba,                         --                    .mem_ba
			mem_ck                   => memory_mem_ck,                         --                    .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                       --                    .mem_ck_n
			mem_cke                  => memory_mem_cke,                        --                    .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                       --                    .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                      --                    .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                      --                    .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                       --                    .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                    --                    .mem_reset_n
			mem_dq                   => memory_mem_dq,                         --                    .mem_dq
			mem_dqs                  => memory_mem_dqs,                        --                    .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                      --                    .mem_dqs_n
			mem_odt                  => memory_mem_odt,                        --                    .mem_odt
			mem_dm                   => memory_mem_dm,                         --                    .mem_dm
			oct_rzqin                => memory_oct_rzqin,                      --                    .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK, --              hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,   --                    .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,   --                    .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,   --                    .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,   --                    .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,   --                    .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,   --                    .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,    --                    .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL, --                    .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL, --                    .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK, --                    .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,   --                    .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,   --                    .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,   --                    .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,     --                    .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,      --                    .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,      --                    .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,     --                    .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,      --                    .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,      --                    .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_hps_io_hps_io_usb1_inst_D0,      --                    .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_hps_io_hps_io_usb1_inst_D1,      --                    .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_hps_io_hps_io_usb1_inst_D2,      --                    .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_hps_io_hps_io_usb1_inst_D3,      --                    .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_hps_io_hps_io_usb1_inst_D4,      --                    .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_hps_io_hps_io_usb1_inst_D5,      --                    .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_hps_io_hps_io_usb1_inst_D6,      --                    .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_hps_io_hps_io_usb1_inst_D7,      --                    .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_hps_io_hps_io_usb1_inst_CLK,     --                    .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_hps_io_hps_io_usb1_inst_STP,     --                    .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_hps_io_hps_io_usb1_inst_DIR,     --                    .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_hps_io_hps_io_usb1_inst_NXT,     --                    .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_0_hps_io_hps_io_spim1_inst_CLK,    --                    .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_hps_io_hps_io_spim1_inst_MOSI,   --                    .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_hps_io_hps_io_spim1_inst_MISO,   --                    .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_hps_io_hps_io_spim1_inst_SS0,    --                    .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,     --                    .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,     --                    .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_hps_io_hps_io_i2c0_inst_SDA,     --                    .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_hps_io_hps_io_i2c0_inst_SCL,     --                    .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_hps_io_hps_io_i2c1_inst_SDA,     --                    .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_hps_io_hps_io_i2c1_inst_SCL,     --                    .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_hps_io_hps_io_gpio_inst_GPIO09,  --                    .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_hps_io_hps_io_gpio_inst_GPIO35,  --                    .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_0_hps_io_hps_io_gpio_inst_GPIO40,  --                    .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_0_hps_io_hps_io_gpio_inst_GPIO53,  --                    .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_hps_io_hps_io_gpio_inst_GPIO54,  --                    .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_hps_io_hps_io_gpio_inst_GPIO61,  --                    .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset_n,               --           h2f_reset.reset_n
			h2f_axi_clk              => clk_clk,                               --       h2f_axi_clock.clk
			h2f_AWID                 => open,                                  --      h2f_axi_master.awid
			h2f_AWADDR               => open,                                  --                    .awaddr
			h2f_AWLEN                => open,                                  --                    .awlen
			h2f_AWSIZE               => open,                                  --                    .awsize
			h2f_AWBURST              => open,                                  --                    .awburst
			h2f_AWLOCK               => open,                                  --                    .awlock
			h2f_AWCACHE              => open,                                  --                    .awcache
			h2f_AWPROT               => open,                                  --                    .awprot
			h2f_AWVALID              => open,                                  --                    .awvalid
			h2f_AWREADY              => open,                                  --                    .awready
			h2f_WID                  => open,                                  --                    .wid
			h2f_WDATA                => open,                                  --                    .wdata
			h2f_WSTRB                => open,                                  --                    .wstrb
			h2f_WLAST                => open,                                  --                    .wlast
			h2f_WVALID               => open,                                  --                    .wvalid
			h2f_WREADY               => open,                                  --                    .wready
			h2f_BID                  => open,                                  --                    .bid
			h2f_BRESP                => open,                                  --                    .bresp
			h2f_BVALID               => open,                                  --                    .bvalid
			h2f_BREADY               => open,                                  --                    .bready
			h2f_ARID                 => open,                                  --                    .arid
			h2f_ARADDR               => open,                                  --                    .araddr
			h2f_ARLEN                => open,                                  --                    .arlen
			h2f_ARSIZE               => open,                                  --                    .arsize
			h2f_ARBURST              => open,                                  --                    .arburst
			h2f_ARLOCK               => open,                                  --                    .arlock
			h2f_ARCACHE              => open,                                  --                    .arcache
			h2f_ARPROT               => open,                                  --                    .arprot
			h2f_ARVALID              => open,                                  --                    .arvalid
			h2f_ARREADY              => open,                                  --                    .arready
			h2f_RID                  => open,                                  --                    .rid
			h2f_RDATA                => open,                                  --                    .rdata
			h2f_RRESP                => open,                                  --                    .rresp
			h2f_RLAST                => open,                                  --                    .rlast
			h2f_RVALID               => open,                                  --                    .rvalid
			h2f_RREADY               => open,                                  --                    .rready
			f2h_axi_clk              => clk_clk,                               --       f2h_axi_clock.clk
			f2h_AWID                 => open,                                  --       f2h_axi_slave.awid
			f2h_AWADDR               => open,                                  --                    .awaddr
			f2h_AWLEN                => open,                                  --                    .awlen
			f2h_AWSIZE               => open,                                  --                    .awsize
			f2h_AWBURST              => open,                                  --                    .awburst
			f2h_AWLOCK               => open,                                  --                    .awlock
			f2h_AWCACHE              => open,                                  --                    .awcache
			f2h_AWPROT               => open,                                  --                    .awprot
			f2h_AWVALID              => open,                                  --                    .awvalid
			f2h_AWREADY              => open,                                  --                    .awready
			f2h_AWUSER               => open,                                  --                    .awuser
			f2h_WID                  => open,                                  --                    .wid
			f2h_WDATA                => open,                                  --                    .wdata
			f2h_WSTRB                => open,                                  --                    .wstrb
			f2h_WLAST                => open,                                  --                    .wlast
			f2h_WVALID               => open,                                  --                    .wvalid
			f2h_WREADY               => open,                                  --                    .wready
			f2h_BID                  => open,                                  --                    .bid
			f2h_BRESP                => open,                                  --                    .bresp
			f2h_BVALID               => open,                                  --                    .bvalid
			f2h_BREADY               => open,                                  --                    .bready
			f2h_ARID                 => open,                                  --                    .arid
			f2h_ARADDR               => open,                                  --                    .araddr
			f2h_ARLEN                => open,                                  --                    .arlen
			f2h_ARSIZE               => open,                                  --                    .arsize
			f2h_ARBURST              => open,                                  --                    .arburst
			f2h_ARLOCK               => open,                                  --                    .arlock
			f2h_ARCACHE              => open,                                  --                    .arcache
			f2h_ARPROT               => open,                                  --                    .arprot
			f2h_ARVALID              => open,                                  --                    .arvalid
			f2h_ARREADY              => open,                                  --                    .arready
			f2h_ARUSER               => open,                                  --                    .aruser
			f2h_RID                  => open,                                  --                    .rid
			f2h_RDATA                => open,                                  --                    .rdata
			f2h_RRESP                => open,                                  --                    .rresp
			f2h_RLAST                => open,                                  --                    .rlast
			f2h_RVALID               => open,                                  --                    .rvalid
			f2h_RREADY               => open,                                  --                    .rready
			h2f_lw_axi_clk           => clk_clk,                               --    h2f_lw_axi_clock.clk
			h2f_lw_AWID              => open,                                  --   h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => open,                                  --                    .awaddr
			h2f_lw_AWLEN             => open,                                  --                    .awlen
			h2f_lw_AWSIZE            => open,                                  --                    .awsize
			h2f_lw_AWBURST           => open,                                  --                    .awburst
			h2f_lw_AWLOCK            => open,                                  --                    .awlock
			h2f_lw_AWCACHE           => open,                                  --                    .awcache
			h2f_lw_AWPROT            => open,                                  --                    .awprot
			h2f_lw_AWVALID           => open,                                  --                    .awvalid
			h2f_lw_AWREADY           => open,                                  --                    .awready
			h2f_lw_WID               => open,                                  --                    .wid
			h2f_lw_WDATA             => open,                                  --                    .wdata
			h2f_lw_WSTRB             => open,                                  --                    .wstrb
			h2f_lw_WLAST             => open,                                  --                    .wlast
			h2f_lw_WVALID            => open,                                  --                    .wvalid
			h2f_lw_WREADY            => open,                                  --                    .wready
			h2f_lw_BID               => open,                                  --                    .bid
			h2f_lw_BRESP             => open,                                  --                    .bresp
			h2f_lw_BVALID            => open,                                  --                    .bvalid
			h2f_lw_BREADY            => open,                                  --                    .bready
			h2f_lw_ARID              => open,                                  --                    .arid
			h2f_lw_ARADDR            => open,                                  --                    .araddr
			h2f_lw_ARLEN             => open,                                  --                    .arlen
			h2f_lw_ARSIZE            => open,                                  --                    .arsize
			h2f_lw_ARBURST           => open,                                  --                    .arburst
			h2f_lw_ARLOCK            => open,                                  --                    .arlock
			h2f_lw_ARCACHE           => open,                                  --                    .arcache
			h2f_lw_ARPROT            => open,                                  --                    .arprot
			h2f_lw_ARVALID           => open,                                  --                    .arvalid
			h2f_lw_ARREADY           => open,                                  --                    .arready
			h2f_lw_RID               => open,                                  --                    .rid
			h2f_lw_RDATA             => open,                                  --                    .rdata
			h2f_lw_RRESP             => open,                                  --                    .rresp
			h2f_lw_RLAST             => open,                                  --                    .rlast
			h2f_lw_RVALID            => open,                                  --                    .rvalid
			h2f_lw_RREADY            => open,                                  --                    .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,                    --            f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq                     --            f2h_irq1.irq
		);

	i2c_opencores_0 : component i2c_opencores
		port map (
			wb_clk_i   => pll_0_outclk0_clk,                                           --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => i2c_0_external_connection_scl_pad_io,                        --           export.export
			sda_pad_io => i2c_0_external_connection_sda_pad_io,                        --                 .export
			wb_adr_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_opencores_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => irq_mapper_002_receiver0_irq                                 -- interrupt_sender.irq
		);

	jtag_uart_nios2 : component Garfield_system_jtag_uart_nios2
		port map (
			clk            => pll_0_outclk0_clk,                                                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                            --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_002_receiver1_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component Garfield_system_nios2_gen2_0
		port map (
			clk                                 => pll_0_outclk0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_nios2 : component Garfield_system_onchip_memory2_nios2
		port map (
			clk        => pll_0_outclk0_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_nios2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_nios2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_nios2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_nios2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_nios2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_nios2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_nios2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                    --       .reset_req
		);

	pll_0 : component Garfield_system_pll_0
		port map (
			refclk   => clk_1_fpga_clock_clk,               --  refclk.clk
			rst      => clk_1_fpga_reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,                  -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	spi_0 : component Garfield_system_spi_0
		port map (
			clk           => pll_0_outclk0_clk,                                        --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_002_receiver3_irq,                             --              irq.irq
			MISO          => spi_0_external_connection_MISO,                           --         external.export
			MOSI          => spi_0_external_connection_MOSI,                           --                 .export
			SCLK          => spi_0_external_connection_SCLK,                           --                 .export
			SS_n          => spi_0_external_connection_SS_n                            --                 .export
		);

	sysid_fpga : component Garfield_system_sysid_fpga
		port map (
			clock    => pll_0_outclk0_clk,                                     --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_fpga_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_fpga_control_slave_address(0)  --              .address
		);

	timer_0_nios2 : component Garfield_system_timer_0_nios2
		port map (
			clk        => pll_0_outclk0_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_timer_0_nios2_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_nios2_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_nios2_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_nios2_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_nios2_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_002_receiver2_irq                        --   irq.irq
		);

	mm_interconnect_0 : component Garfield_system_mm_interconnect_0
		port map (
			pll_0_outclk0_clk                              => pll_0_outclk0_clk,                                               --                            pll_0_outclk0.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                  -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                                --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                            --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                             --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                                   --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                               --                                         .readdata
			nios2_gen2_0_data_master_readdatavalid         => nios2_gen2_0_data_master_readdatavalid,                          --                                         .readdatavalid
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                                  --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                              --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                            --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                         --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                     --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                            --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                        --                                         .readdata
			nios2_gen2_0_instruction_master_readdatavalid  => nios2_gen2_0_instruction_master_readdatavalid,                   --                                         .readdatavalid
			Garfield_GPIO_s1_address                       => mm_interconnect_0_garfield_gpio_s1_address,                      --                         Garfield_GPIO_s1.address
			Garfield_GPIO_s1_write                         => mm_interconnect_0_garfield_gpio_s1_write,                        --                                         .write
			Garfield_GPIO_s1_readdata                      => mm_interconnect_0_garfield_gpio_s1_readdata,                     --                                         .readdata
			Garfield_GPIO_s1_writedata                     => mm_interconnect_0_garfield_gpio_s1_writedata,                    --                                         .writedata
			Garfield_GPIO_s1_chipselect                    => mm_interconnect_0_garfield_gpio_s1_chipselect,                   --                                         .chipselect
			Garfield_lighting_s1_address                   => mm_interconnect_0_garfield_lighting_s1_address,                  --                     Garfield_lighting_s1.address
			Garfield_lighting_s1_write                     => mm_interconnect_0_garfield_lighting_s1_write,                    --                                         .write
			Garfield_lighting_s1_readdata                  => mm_interconnect_0_garfield_lighting_s1_readdata,                 --                                         .readdata
			Garfield_lighting_s1_writedata                 => mm_interconnect_0_garfield_lighting_s1_writedata,                --                                         .writedata
			Garfield_lighting_s1_chipselect                => mm_interconnect_0_garfield_lighting_s1_chipselect,               --                                         .chipselect
			i2c_opencores_0_avalon_slave_0_address         => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,        --           i2c_opencores_0_avalon_slave_0.address
			i2c_opencores_0_avalon_slave_0_write           => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,          --                                         .write
			i2c_opencores_0_avalon_slave_0_readdata        => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,       --                                         .readdata
			i2c_opencores_0_avalon_slave_0_writedata       => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,      --                                         .writedata
			i2c_opencores_0_avalon_slave_0_waitrequest     => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv,            --                                         .waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect      => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect,     --                                         .chipselect
			jtag_uart_nios2_avalon_jtag_slave_address      => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_address,     --        jtag_uart_nios2_avalon_jtag_slave.address
			jtag_uart_nios2_avalon_jtag_slave_write        => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_nios2_avalon_jtag_slave_read         => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_nios2_avalon_jtag_slave_readdata     => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_nios2_avalon_jtag_slave_writedata    => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_nios2_avalon_jtag_slave_waitrequest  => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_nios2_avalon_jtag_slave_chipselect   => mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_chipselect,  --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,          --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,            --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,             --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,         --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,        --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,       --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,      --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,      --                                         .debugaccess
			Onboard_Button_s1_address                      => mm_interconnect_0_onboard_button_s1_address,                     --                        Onboard_Button_s1.address
			Onboard_Button_s1_write                        => mm_interconnect_0_onboard_button_s1_write,                       --                                         .write
			Onboard_Button_s1_readdata                     => mm_interconnect_0_onboard_button_s1_readdata,                    --                                         .readdata
			Onboard_Button_s1_writedata                    => mm_interconnect_0_onboard_button_s1_writedata,                   --                                         .writedata
			Onboard_Button_s1_chipselect                   => mm_interconnect_0_onboard_button_s1_chipselect,                  --                                         .chipselect
			Onboard_DipSW_s1_address                       => mm_interconnect_0_onboard_dipsw_s1_address,                      --                         Onboard_DipSW_s1.address
			Onboard_DipSW_s1_write                         => mm_interconnect_0_onboard_dipsw_s1_write,                        --                                         .write
			Onboard_DipSW_s1_readdata                      => mm_interconnect_0_onboard_dipsw_s1_readdata,                     --                                         .readdata
			Onboard_DipSW_s1_writedata                     => mm_interconnect_0_onboard_dipsw_s1_writedata,                    --                                         .writedata
			Onboard_DipSW_s1_chipselect                    => mm_interconnect_0_onboard_dipsw_s1_chipselect,                   --                                         .chipselect
			Onboard_LED_s1_address                         => mm_interconnect_0_onboard_led_s1_address,                        --                           Onboard_LED_s1.address
			Onboard_LED_s1_write                           => mm_interconnect_0_onboard_led_s1_write,                          --                                         .write
			Onboard_LED_s1_readdata                        => mm_interconnect_0_onboard_led_s1_readdata,                       --                                         .readdata
			Onboard_LED_s1_writedata                       => mm_interconnect_0_onboard_led_s1_writedata,                      --                                         .writedata
			Onboard_LED_s1_chipselect                      => mm_interconnect_0_onboard_led_s1_chipselect,                     --                                         .chipselect
			onchip_memory2_nios2_s1_address                => mm_interconnect_0_onchip_memory2_nios2_s1_address,               --                  onchip_memory2_nios2_s1.address
			onchip_memory2_nios2_s1_write                  => mm_interconnect_0_onchip_memory2_nios2_s1_write,                 --                                         .write
			onchip_memory2_nios2_s1_readdata               => mm_interconnect_0_onchip_memory2_nios2_s1_readdata,              --                                         .readdata
			onchip_memory2_nios2_s1_writedata              => mm_interconnect_0_onchip_memory2_nios2_s1_writedata,             --                                         .writedata
			onchip_memory2_nios2_s1_byteenable             => mm_interconnect_0_onchip_memory2_nios2_s1_byteenable,            --                                         .byteenable
			onchip_memory2_nios2_s1_chipselect             => mm_interconnect_0_onchip_memory2_nios2_s1_chipselect,            --                                         .chipselect
			onchip_memory2_nios2_s1_clken                  => mm_interconnect_0_onchip_memory2_nios2_s1_clken,                 --                                         .clken
			spi_0_spi_control_port_address                 => mm_interconnect_0_spi_0_spi_control_port_address,                --                   spi_0_spi_control_port.address
			spi_0_spi_control_port_write                   => mm_interconnect_0_spi_0_spi_control_port_write,                  --                                         .write
			spi_0_spi_control_port_read                    => mm_interconnect_0_spi_0_spi_control_port_read,                   --                                         .read
			spi_0_spi_control_port_readdata                => mm_interconnect_0_spi_0_spi_control_port_readdata,               --                                         .readdata
			spi_0_spi_control_port_writedata               => mm_interconnect_0_spi_0_spi_control_port_writedata,              --                                         .writedata
			spi_0_spi_control_port_chipselect              => mm_interconnect_0_spi_0_spi_control_port_chipselect,             --                                         .chipselect
			sysid_fpga_control_slave_address               => mm_interconnect_0_sysid_fpga_control_slave_address,              --                 sysid_fpga_control_slave.address
			sysid_fpga_control_slave_readdata              => mm_interconnect_0_sysid_fpga_control_slave_readdata,             --                                         .readdata
			timer_0_nios2_s1_address                       => mm_interconnect_0_timer_0_nios2_s1_address,                      --                         timer_0_nios2_s1.address
			timer_0_nios2_s1_write                         => mm_interconnect_0_timer_0_nios2_s1_write,                        --                                         .write
			timer_0_nios2_s1_readdata                      => mm_interconnect_0_timer_0_nios2_s1_readdata,                     --                                         .readdata
			timer_0_nios2_s1_writedata                     => mm_interconnect_0_timer_0_nios2_s1_writedata,                    --                                         .writedata
			timer_0_nios2_s1_chipselect                    => mm_interconnect_0_timer_0_nios2_s1_chipselect                    --                                         .chipselect
		);

	irq_mapper : component Garfield_system_irq_mapper
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq0_irq  --    sender.irq
		);

	irq_mapper_001 : component Garfield_system_irq_mapper
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	irq_mapper_002 : component Garfield_system_irq_mapper_002
		port map (
			clk           => pll_0_outclk0_clk,              --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_002_receiver0_irq,   -- receiver0.irq
			receiver1_irq => irq_mapper_002_receiver1_irq,   -- receiver1.irq
			receiver2_irq => irq_mapper_002_receiver2_irq,   -- receiver2.irq
			receiver3_irq => irq_mapper_002_receiver3_irq,   -- receiver3.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_1_fpga_reset_reset_n_ports_inv, -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	clk_1_fpga_reset_reset_n_ports_inv <= not clk_1_fpga_reset_reset_n;

	mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_nios2_avalon_jtag_slave_write;

	mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv <= not i2c_opencores_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_onboard_led_s1_write_ports_inv <= not mm_interconnect_0_onboard_led_s1_write;

	mm_interconnect_0_onboard_button_s1_write_ports_inv <= not mm_interconnect_0_onboard_button_s1_write;

	mm_interconnect_0_onboard_dipsw_s1_write_ports_inv <= not mm_interconnect_0_onboard_dipsw_s1_write;

	mm_interconnect_0_timer_0_nios2_s1_write_ports_inv <= not mm_interconnect_0_timer_0_nios2_s1_write;

	mm_interconnect_0_garfield_lighting_s1_write_ports_inv <= not mm_interconnect_0_garfield_lighting_s1_write;

	mm_interconnect_0_garfield_gpio_s1_write_ports_inv <= not mm_interconnect_0_garfield_gpio_s1_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Garfield_system
